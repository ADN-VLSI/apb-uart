module apb_uart_tb;

  initial begin
    $display("This is a placeholder testbench for apb_uart.");
    $finish;
  end

endmodule
